*  Generated for: PrimeSim
*  Design library name: CSA
*  Design cell name: test_8bit_CSA
*  Design view name: schematic
.lib 'saed32nm.lib' TT

*Custom Compiler Version S-2021.09
*Fri Feb 25 20:05:21 2022

.global gnd!
********************************************************************************
* Library          : CSA
* Cell             : inverter
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt inverter in out vdc gnd_1
xm0 out in gnd_1 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm1 out in vdc vdc p105 w=0.1u l=0.03u nf=1 m=1
.ends inverter

********************************************************************************
* Library          : CSA
* Cell             : FA
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt fa a b carry cin gnd_1 sum vdc1 vdc2
xi7 net75 net67 vdc2 gnd_1 inverter
xi6 cin net52 vdc2 gnd_1 inverter
xi1 b net24 vdc1 gnd_1 inverter
xi0 a net22 vdc1 gnd_1 inverter
xm14 b net67 carry gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm13 cin net75 carry gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm9 net52 net75 sum gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm12 cin net67 sum gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm3 net24 a net75 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm2 b net22 net75 gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm16 b net75 carry vdc2 p105 w=0.1u l=0.03u nf=1 m=1
xm15 cin net67 carry vdc2 p105 w=0.1u l=0.03u nf=1 m=1
xm11 net52 net67 sum vdc2 p105 w=0.1u l=0.03u nf=1 m=1
xm10 cin net75 sum vdc2 p105 w=0.1u l=0.03u nf=1 m=1
xm5 net24 net22 net75 vdc1 p105 w=0.1u l=0.03u nf=1 m=1
xm4 b a net75 vdc1 p105 w=0.1u l=0.03u nf=1 m=1
.ends fa

********************************************************************************
* Library          : CSA
* Cell             : 4bit_RCA
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt _4bit_rca a0 a1 a2 a3 b0 b1 b2 b3 cin cout gnd_1 s0 s1 s2 s3 vdc
xi3 a3 b3 cout net25 gnd_1 s3 vdc vdc fa
xi2 a2 b2 net25 net17 gnd_1 s2 vdc vdc fa
xi1 a1 b1 net17 net9 gnd_1 s1 vdc vdc fa
xi0 a0 b0 net9 cin gnd_1 s0 vdc vdc fa
.ends _4bit_rca

********************************************************************************
* Library          : CSA
* Cell             : XOR
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt xor a b gnd_1 out vdc
xm1 a net10 out gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm0 net12 b out gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm3 a b out vdc p105 w=0.1u l=0.03u nf=1 m=1
xm2 net12 net10 out vdc p105 w=0.1u l=0.03u nf=1 m=1
xi5 b net10 vdc gnd_1 inverter
xi4 a net12 vdc gnd_1 inverter
.ends xor

********************************************************************************
* Library          : CSA
* Cell             : 2_input_AND
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt _2_input_and a b gnd_1 out vdc
xi5 b net18 vdc gnd_1 inverter
xm3 out b a gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm4 out net18 b gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
.ends _2_input_and

********************************************************************************
* Library          : CSA
* Cell             : BtoE1
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt btoe1 p0 p1 p2 p3 q0 q1 q2 q3 qcout vdc gnd_1
xi0 p0 q0 vdc gnd_1 inverter
xi3 net33 p3 gnd_1 q3 vdc xor
xi2 p0 p1 gnd_1 q1 vdc xor
xi1 net28 p2 gnd_1 q2 vdc xor
xi6 net33 p3 gnd_1 qcout vdc _2_input_and
xi5 net28 p2 gnd_1 net33 vdc _2_input_and
xi4 p0 p1 gnd_1 net28 vdc _2_input_and
.ends btoe1

********************************************************************************
* Library          : CSA
* Cell             : 2:1_MUX
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt _2:1_mux in1 in2 out signal vdc gnd_1
xm1 in2 signal out gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm0 in1 net10 out gnd_1 n105 w=0.1u l=0.03u nf=1 m=1
xm3 in1 signal out vdc p105 w=0.1u l=0.03u nf=1 m=1
xm2 in2 net10 out net24 p105 w=0.1u l=0.03u nf=1 m=1
xi4 signal net10 vdc gnd_1 inverter
.ends _2:1_mux

********************************************************************************
* Library          : CSA
* Cell             : 2:1_mux_array
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt _2:1_mux_array cout q4 q5 q6 q7 qcout s4 s5 s6 s7 slc_signal z4 z5 z6 z7
+  zcout gnd_1 vdc
xi4 zcout qcout cout slc_signal vdc gnd_1 _2:1_mux
xi3 z4 q4 s4 slc_signal vdc gnd_1 _2:1_mux
xi2 z7 q7 s7 slc_signal vdc gnd_1 _2:1_mux
xi1 z6 q6 s6 slc_signal vdc gnd_1 _2:1_mux
xi0 z5 q5 s5 slc_signal vdc gnd_1 _2:1_mux
.ends _2:1_mux_array

********************************************************************************
* Library          : CSA
* Cell             : 8_bit_CSAwithBtoE1converter
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt _8_bit_csawithbtoe1converter a0 a1 a2 a3 a4 a5 a6 a7 b0 b1 b2 b3 b4 b5
+ b6 b7 cout gnd_1 s0 s1 s2 s3 s4 s5 s6 s7 vdc
xi1 a4 a5 a6 a7 b4 b5 b6 b7 gnd_1 net51 gnd_1 net45 net46 net47 net49 vdc
+ _4bit_rca
xi0 a0 a1 a2 a3 b0 b1 b2 b3 gnd_1 net43 gnd_1 s0 s1 s2 s3 vdc _4bit_rca
xi2 net45 net46 net47 net49 net53 net55 net57 net58 net61 vdc gnd_1 btoe1
xi3 cout net53 net55 net57 net58 net61 s4 s5 s6 s7 net43 net45 net46 net47 net49
+ net51 gnd_1 vdc _2:1_mux_array
.ends _8_bit_csawithbtoe1converter

********************************************************************************
* Library          : CSA
* Cell             : test_8bit_CSA
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
xi0 a0 a1 a2 a3 a4 a5 a6 a7 b0 b1 b2 b3 b4 b5 b6 b7 cout gnd! s0 s1 s2 s3 s4 s5
+ s6 s7 net29 _8_bit_csawithbtoe1converter
v2 net29 gnd! dc=.8
v18 b7 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 256u 512u )
v17 b0 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 2u 4u )
v16 b1 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 4 8 )
v15 b2 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 8u 16u )
v14 b3 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 16u 32u )
v13 b4 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 32u 64u )
v12 b5 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 64u 128u )
v11 b6 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 128u 256u )
v10 a0 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 1.5u 3u )
v9 a7 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 192u 384u )
v8 a6 gnd! dc=0 pulse ( 1.2 0 0 0.1u .1u 96u 192u )
v7 a5 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 48u 96u )
v6 a4 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 24u 48u )
v5 a3 gnd! dc=0 pulse ( 1.2 0 0 .1u .1u 12u 24u )
v4 a2 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 6u 12u )
v3 a1 gnd! dc=0 pulse ( 1.20 0 0 .1u .1u 3u 6u )








.tran '1u' '500u' name=tran

.option primesim_remove_probe_prefix = 0
.probe v(*) i(*) level=1
.probe tran v(a0) v(a1) v(a2) v(a3) v(a4) v(a5) v(a6) v(a7) v(b0) v(b1) v(b2)
+ v(b3) v(b4) v(b5) v(b6) v(b7) v(cout) v(s0) v(s1) v(s2) v(s3) v(s4) v(s5)
+ v(s6) v(s7)

.temp 25



.option primesim_output=wdf


.option parhier = LOCAL






.end
