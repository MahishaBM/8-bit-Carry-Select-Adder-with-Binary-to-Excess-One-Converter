*  Generated for: PrimeSim
*  Design library name: CSA
*  Design cell name: test_inverter
*  Design view name: schematic
.lib 'saed32nm.lib' TT

*Custom Compiler Version S-2021.09
*Sun Feb 20 15:02:48 2022

.global gnd!
********************************************************************************
* Library          : CSA
* Cell             : inverter
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
.subckt inverter net3 net7 net8 net9
xm0 net7 net8 net3 net3 n105 w=0.1u l=0.03u nf=1 m=1
xm1 net7 net8 net9 net9 p105 w=0.1u l=0.03u nf=1 m=1
.ends inverter

********************************************************************************
* Library          : CSA
* Cell             : test_inverter
* View             : schematic
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
xi0 gnd! out in net5 inverter
v2 net5 gnd! dc=1.2
v3 in gnd! dc=0 pulse ( 0 1.05 0 0.1u 0.1u 10u 20u )








.tran '1u' '20u' name=tran

.option primesim_remove_probe_prefix = 0
.probe v(*) i(*) level=1
.probe tran v(in) v(out)

.temp 25



.option primesim_output=wdf


.option parhier = LOCAL






.end
